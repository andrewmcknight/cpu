// shift_left_2: Logical left shift by 2 bits for 32-bit inputs. Inputs: in. Outputs: out.

module shift_left_2(out, in);
    input [31:0] in;
    output [31:0] out;

    assign out = {in[29:0], 2'b00};
endmodule
